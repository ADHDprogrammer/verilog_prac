module moduleName (
    // no input
    );

    
    
endmodule